-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Nov  2 16:22:44 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maq_estados IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        LED3 : OUT STD_LOGIC;
        LED2 : OUT STD_LOGIC;
        LED1 : OUT STD_LOGIC;
        LED0 : OUT STD_LOGIC
    );
END maq_estados;

ARCHITECTURE BEHAVIOR OF maq_estados IS
    TYPE type_fstate IS (A,B,C,D,E,F,G);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            LED3 <= '0';
            LED2 <= '0';
            LED1 <= '0';
            LED0 <= '0';
        ELSE
            LED3 <= '0';
            LED2 <= '0';
            LED1 <= '0';
            LED0 <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((x = '0')) THEN
                        reg_fstate <= B;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= E;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    LED3 <= '0';

                    LED2 <= '0';

                    LED0 <= '0';

                    LED1 <= '0';
                WHEN B =>
                    reg_fstate <= C;

                    LED3 <= '0';

                    LED2 <= '1';

                    LED0 <= '0';

                    LED1 <= '1';
                WHEN C =>
                    IF ((x = '0')) THEN
                        reg_fstate <= D;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= G;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C;
                    END IF;

                    LED3 <= '1';

                    LED2 <= '1';

                    LED0 <= '1';

                    LED1 <= '1';
                WHEN D =>
                    reg_fstate <= A;

                    LED3 <= '1';

                    LED2 <= '0';

                    LED0 <= '1';

                    LED1 <= '0';
                WHEN E =>
                    reg_fstate <= F;

                    LED3 <= '1';

                    LED2 <= '0';

                    LED0 <= '0';

                    LED1 <= '0';
                WHEN F =>
                    reg_fstate <= C;

                    LED3 <= '1';

                    LED2 <= '1';

                    LED0 <= '0';

                    LED1 <= '0';
                WHEN G =>
                    reg_fstate <= A;

                    LED3 <= '1';

                    LED2 <= '1';

                    LED0 <= '0';

                    LED1 <= '1';
                WHEN OTHERS => 
                    LED3 <= 'X';
                    LED2 <= 'X';
                    LED1 <= 'X';
                    LED0 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
